library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity T13_ConcurrentStatement is
end entity;

architecture sim of T13_ConcurrentStatement is
	signal Uns : unsigned(5 downto 0):=(others=>'0');
	signal Mul1: unsigned(7 downto 0);
	signal Mul2: unsigned(7 downto 0);
	
begin

	process is
	begin
		Uns <= Uns +1;
		wait on Uns;
		
	    
	end process;
	process(Uns) is 
	begin
		Mul1 <= Uns & "00";
		
	end process;	
	Mul2 <= Uns & "00";
end architecture;